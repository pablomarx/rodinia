module top;

	wire clk;
	(* BEL="IOTILE(04,09):alta_rio00", keep *) /* PIN_46 */
	GENERIC_IOB #(.INPUT_USED(1), .OUTPUT_USED(0)) clk_ibuf (.O(clk));

	wire [7:0] leds;
	(* BEL="IOTILE(02,01):alta_rio02", keep *)	/* PIN_11 */
	GENERIC_IOB #(.INPUT_USED(0), .OUTPUT_USED(1)) led7_obuf (.I(leds[7]));
	(* BEL="IOTILE(07,01):alta_rio00", keep *)	/* PIN_09 */
	GENERIC_IOB #(.INPUT_USED(0), .OUTPUT_USED(1)) led6_obuf (.I(leds[6]));
	(* BEL="IOTILE(06,09):alta_rio02", keep *)  /* PIN_06 */
	GENERIC_IOB #(.INPUT_USED(0), .OUTPUT_USED(1)) led5_obuf (.I(leds[5]));
	(* BEL="IOTILE(01,09):alta_rio01", keep *)  /* PIN_05 */
	GENERIC_IOB #(.INPUT_USED(0), .OUTPUT_USED(1)) led4_obuf (.I(leds[4]));
	(* BEL="IOTILE(00,09):alta_rio00", keep *)	/* PIN_04 */
	GENERIC_IOB #(.INPUT_USED(0), .OUTPUT_USED(1)) led3_obuf (.I(leds[3]));
	(* BEL="IOTILE(00,09):alta_rio02", keep *)	/* PIN_03 */
	GENERIC_IOB #(.INPUT_USED(0), .OUTPUT_USED(1)) led2_obuf (.I(leds[2]));
	(* BEL="IOTILE(01,09):alta_rio03", keep *)	/* PIN_02 */
	GENERIC_IOB #(.INPUT_USED(0), .OUTPUT_USED(1)) led1_obuf (.I(leds[1]));
	(* BEL="IOTILE(02,09):alta_rio00", keep *)	/* PIN_01 */
	GENERIC_IOB #(.INPUT_USED(0), .OUTPUT_USED(1)) led0_obuf (.I(leds[0]));

reg [25:0] ctr;
always @(posedge clk)
	ctr <= ctr + 1'b1;

//assign leds = ctr[25:18];

GENERIC_BRAM ram_inst(
	.AddressA(ctr[24:13]),
	.DataOutA(leds),
	.WeRenA(1'b0),
	.AsyncReset0(1'b0),
	.Clk0(clk),
);

defparam ram_inst.INIT_VAL = 4608'b011011101001001110111111001111001001101111111000011010000010101010010011110100100101011101000011100001001000111010101101100101110100000010111000111100010111101011000000000101001111101110011110110101001110001101100011111110110001101001001110011001000010011001010110101100011000001011001011001011100001000100100000001101011110000110010011010000101001001111001100110000000101110111001111101010010001001010010110010100011001001101000100000110001100011101011110010000010100111110111011000000010110001000000001100001101011000010000011010110011101011110110000110100001100100001010101100110110111010001110000100110100011011101010110011000111111001010110010011110010111101010000000001100011010110001110000111011111110101110100010000101011010111100100111111100100010010111100000001001010011100100101111110000010011100110101001111101000011100110101100100000111101100100010111001011110010010100101101010110000101111111001111000010100101011011010001110111110000101011100111010001110111111111110001010011100011100111001010001110110010000101111101000010100101101110011010001101101000111100111011101001011110011011011111010011111100111001110111101100010000111100000110000010001101011010001011110001100011011101010011001011011111000010000000111001111100100101101001010100101100001100111010000110010001101101110111011000010111000000010110001110101110110111001010000001100011110000111010010111001011100000111110110011100011011110011101111101101000111001110111100110010000111111010000010001111000101010101101110001001011101001000101101111001000001001000010001000000110111110111101011010011011110000011011000101101101111000001111010001011010010111101000011011000111100001001100101100110101110001001101101000010110000011111000001011101100111101101101010101100000011100000111111000011100001011010011011101100010011001010011101000110000100001001111001010000000100010111110111111101000010101011110101111011111010001001101010101101011010001111010000001100111110011111000100111001001000000001000100000001101110111010011001001010010100110111010011100101001101011101000010011110011011011101101010001110011110101110011101101001111111000110110110100010111111110101110000111100110100100001001001000000011001000110100101111001111000111010111100011000011100011101000110011000010100101110000011100110110000101001100111000001010101101101110011000101110110100001001011000101011010101001101111100100111001110000010011010101010100100101110000111110111000010010111110011011001011001100000010011011111100010011100011101110100000110011101100111111110011111010011111011101011011001001110110000010100100001100111101110100000110001011111000010011011110100010011111111010000101010101110111010010101100001011010001001010001110001100010001000111101000011110001100011011101111011001001001110011010001100001101110010111100011000001011100011011010101001101001110100011110110010110101100010101011001001000000110011101011100010011110111110001101000000011100001001110100100111101011000010100011011001010011010010101100101000010011010111110001110000110010100111001001011011100010101010000101001101000110110101110100010111000010011100111101100100010110001110011011001100100000010011011101010110111111010000101010000011111101001000010011010010000111010000100011111111001111100000100110011000001011000100001111000110110010001001101000000110101011011011110100001110100111100010100100110000010001001100011101110100110011111101010010001101110100101101011011010000101001011010010011011011001110101111011111011100010010010111100101111111101110110001010101110100101000010111100011110110111001011100111111110011100100001010010011011011100100111010001000111010111100001010001000011100010011010100000110001100101100100010000111111000111010011100111011100111000010110000110110101011101001011101111101000010001011011100011100011111110010101110010101000010010110000111100001001100010111100111011011001110001101000000001010011100000001010100010000011011111011010011000010111100110111000011100111110111010101010000000010010011110100011111011011011100010011011100001110110111000101010001101101110100000000111110100100001111000110101111100010100011101000111011011001110010100100110001011101010100110000001000010111110101000101000110101100100010101001000111100101100100110000001111011100110001101010101110110101111001100001001101011100000011001111011100111011001101000000000010111011011000111101011101111111100011111111000111001100010001000000110110111010000001001011010110011110010010110101011100100101101001011000111110111100001101111110000110011100110110001000011101000100111000100111001001010110100101011101010101111000001000100010100000110000000110111000110000010000011101000011;


endmodule
