module top;

	wire clk;
	(* BEL="IOTILE(40,12):alta_rio02", keep *) /* PIN_112 */
	GENERIC_IOB #(.INPUT_USED(1), .OUTPUT_USED(0)) clk_ibuf (.O(clk));

	wire [7:0] leds;
	(* BEL="IOTILE(38,00):alta_rio03", keep *)	/* PIN_87 */
	GENERIC_IOB #(.INPUT_USED(0), .OUTPUT_USED(1)) led7_obuf (.I(leds[7]));
	(* BEL="IOTILE(38,00):alta_rio02", keep *)	/* PIN_88 */
	GENERIC_IOB #(.INPUT_USED(0), .OUTPUT_USED(1)) led6_obuf (.I(leds[6]));
	(* BEL="IOTILE(40,02):alta_rio01", keep *)  /* PIN_89 */
	GENERIC_IOB #(.INPUT_USED(0), .OUTPUT_USED(1)) led5_obuf (.I(leds[5]));
	(* BEL="IOTILE(40,02):alta_rio00", keep *)  /* PIN_90 */
	GENERIC_IOB #(.INPUT_USED(0), .OUTPUT_USED(1)) led4_obuf (.I(leds[4]));
	(* BEL="IOTILE(40,03):alta_rio01", keep *)	/* PIN_91 */
	GENERIC_IOB #(.INPUT_USED(0), .OUTPUT_USED(1)) led3_obuf (.I(leds[3]));
	(* BEL="IOTILE(40,03):alta_rio00", keep *)	/* PIN_92 */
	GENERIC_IOB #(.INPUT_USED(0), .OUTPUT_USED(1)) led2_obuf (.I(leds[2]));
	(* BEL="IOTILE(40,04):alta_rio01", keep *)	/* PIN_93 */
	GENERIC_IOB #(.INPUT_USED(0), .OUTPUT_USED(1)) led1_obuf (.I(leds[1]));
	(* BEL="IOTILE(40,04):alta_rio00", keep *)	/* PIN_94 */
	GENERIC_IOB #(.INPUT_USED(0), .OUTPUT_USED(1)) led0_obuf (.I(leds[0]));

reg [25:0] ctr;
always @(posedge clk)
	ctr <= ctr + 1'b1;

//assign leds = ctr[25:18];

alta_bram9k ram_inst(
	.AddressA(ctr[24:13]),
	.DataOutA(leds),
	.WeA(1'b0),
	.ReA(1'b1),
	.AsyncReset0(1'b0),
	.Clk0(clk),
	.ClkEn0(1'b1),
);

defparam ram_inst.INIT_VAL = 9216'h4d8c09c2f983e412ebf7a005a4f86a6dd527348fd73608837aabf94f06cfdbab1f702c5796451a35f4cc21049420ac6c21512d9d1ea94bcc8cc5b4a47ae75f35764ff05676323ee1de6ad0e18ac7c494b1dc5899d6e619bfaff03fe1949f154a7bcb4bd955a7fde964d841ef35fc6830c5d496f96f15e9ad03645be351cb300cbb14e130a65db0fb0bb9c711712a8c84e7eea0a2c7461e7ae7ad02f5464894d6798e41514a9a87b1912af07f49b215bd150f5d495e2eb1793f974dd265ca0be094cebcb3c2c2e099aed8b38e344e9335fb8c41111a7d45dbf3c456e7a867372685291033e68db115dc197e510e92f7195780c790d5defefde00338a097ae2ee8b9ab2b3cd453082350cb6e28b59066af594cbb68ffa421b657ee89b5e5057c84c1507fe0591ec592e95e77a9d4f653cc3dbca25258cdc46cbec21809a2d68febc93b6d9629d766ac7043cb737979913f34f6a774d2d3262c32d8e6c7c5cc315ed02503638826e997d42580c16638b1eacbb2977cc6a735bd67ba99d9f474e08751d9ae2e4eb6283e68793f9aa9ed9a933121b985167038bddfb892b2c63ccb03471a4ddf43f1c82813da80c687434731fb9de631e9c5b6e29acfea466605057700df86663373320e40b41d8410879d0132820602bda0ad3668b7709369782af9090d6d86c168470db32546b186783d14cdd7a3aaac1c1d352248e7e167cdbec13977423c53491ee497e2a85acb6a259e00e077957242dcad6850319b410370fd88783f4030e45b51b520674d56d2eae66ef38eb8857ef1ccae170fecc1ac72fb0d8115168d529ea7ae5cad90929c54b7118172a673d685059257424ac14813f40e3c4fe8ee0464b072309a402a1fc0da24fcc264d4cf9ea0e21d7bdc57b712b695a787fe0d2a47387bb911c453680377fb990208215c017451f18ec65436bd8963b6d3e496e2ba055fd307dcec4afcb50175b39267da2c4fedbe969e23a2f200bb1e5b94ddf738d5725df08c2fc2baa0dac187c54b8e2ec74d8ad2f26c22499a8a5111af06067269e25c72234fdccc0ee1115e61b1f07365bb3a8ca8763b85e986fe179c4033853410ba8695371dff4c75773a966cb7d045b7fa56d6446aa2244f552e13de484a118ea0f579efde2fb4b9d9f85d43a54a560979c8a02d25717b3cad09c5525bc18667c0dc56c7e7c8a677dfbcbdbe12201e5562793116f369b37a8f6dcc67e10a7d55f39fce24663de222bdb687fc6b0be2e5c54c471df0c3ae18851967a330bd40efb23af58ffc04dba93a32d4149250a71818cdeeb8b95a98f2c7de0ee1fe77a4d818cdc26d134c4b0ca2fda4f35ecb0991897f25de6ad582a5bdf7d64da193a62e75f0cf95ece3a5b81d7db8167955b33475636728bd29ab95da4da1c614256fbbcacc245e31fdff1005266eaf5dee25d29350500ab7e3c7105ff4c5170cf4905e7bab3186b47cdd1ff2401ec87aa3f72cfb68c8c8e2d0bd9b83b6b4f724b37ae1558cc63777bd0f6f75ac71f6ed7dd17aa4acc3c7b63513fc1356359dad4e453c04dbddb5076c6b20282270507accb0030dc8284136010f8911ea0f26ab93a12e737285a8daa32aeb9c177f5192465b0e48e5efb15089da;


endmodule
