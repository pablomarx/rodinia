`timescale 1ns/1ps
module prom(
   input clka,
   input clkb,

   input [12:0] addra,
   input [12:0] addrb,

   output [35:0] douta,
   output [35:0] doutb,

   input wea,
   input [35:0] dina
);


alta_bram9k ram_inst(
.DataOutA(douta), .DataInA(dina), .AddressA(addra), .ByteEnA(1'b0), .Clk0(clka), .ClkEn0(1'b1),
.AsyncReset0(1'b0), .AddressStallA(1'b0), .WeA(wea), .ReA(1'b1),

.DataOutB(doutb), .DataInB(), .AddressB(addrb), .ByteEnB(1'b0), .Clk1(clkb), .ClkEn1(1'b1),
.AsyncReset1(1'b0), .AddressStallB(1'b0), .WeB(1'b0), .ReB(1'b1),
);

defparam ram_inst.INIT_VAL = 9216'h86d8c5636b2e163e62b874a187cb29c76ac21448535bc5f2f9185fa192c20fcded0552b1f7510ece6fd171b31df39371f41d3a1c50c38c187edb591401ba60d532c6f862894575941e1bd0a85043d45bbdd08b7f63d6e13f3687ca69612028fee4fd2d6969f3cb67c6bcac9be184a1e666a7c5b70b830d38ca54b1f75da1170bc54e731170ad561c9e24fe778e281040dba9f97f3bb4b27979a00f611a7257acf506bc8e92299328a72784a2000e875c0f29b6d07dd8cf631f0e30b5dbf052d1409868ede69c00aa0731852a2ccf6ef133b993ec74b8f206a945ef617adb3fec5fa4b9d97ac4541ef6b68815270136a61d0e86cfd08588a95ddcc29c2c99413bd85990d42bf63863875a01c6d2501e147d6e18dc5a9cc5388363a3450be9fcc7f4cab46e4e7dde884ed9765e8a052e71ff70c8db6f6ead537ffa43ff939cab1988956ea5da06864c6541d2ba5642da988bd69b8cd7db6cdd0b91422880b9771740498cbc84e5ddfce8dd6e4045b1e2ec1e97421657408bb6829ed401bf9136b74c850cbd5ebdffa953e4ffba354eccce7da84f8239636ee0a4a32f332c4e33943a0cfdb200f907269f91e80f2d06761bacb9c21d91248b1d0b5bca4d9e62f15e0a26c807b385c1ff5cd0333475bc6fcbc531647a3c396958bd51ed36ebc10bbcf86ce22de163ae064d39ada69ea8d1dae334033d26db14e834ffacc1441b0006cdbbcdc57b82de5d8218e75a7d776ca21c0fc21270008b8b7cd9d80c220bbaff424e253be7a13756c5c5f773609ee34ff3ef792dc4989b5309e02ae375a86f8db8fca8229bc3c2ba6ddf4e108e37cd53764bc98f39b796a8294abed665edc9773b4ddab91637a0ae57f9ec87659aac0feb0987a5d08e47f302ac040dfaec405df83c6d69c532a98e67bcaf6ee923a84c4c968617ca772184afc4a37cb996812371d0cd92b7555154d1aa4e45db2f0d7113a4ab18a5e7b93963396c2089554244d20d2e9c84bb410143a8329008efe544acbd4379bd3b31597e747bcf71ab0fe0da7bd344dbd160e4f6cc88fd774165ff41415bd92bf18f11ffb6a75d7b9dfc1ec7e6dc8cf63b1348e861a22a3184c3c07ed8292be445c59ac315ed6ea9795fed300dd58cf406c500d58776d189a483282d2f4d31ca39e250cc228c264f120a9f905273bdfa0b56f34ce26f5a72544584d85459f7944b6f61e179daadb56d5f1a9ad7ba612739e8d0c95e7f3c1a7809c7eca428a99f866ec2759a9644adc8e629f37a91adbd3ab586dfb0ee9d2eee13807f925194278aa27d0d1b894ac85393ca8de2d7bc8444a87dacc37332eb3bce4889f94df80a5cbc015402c466fc811b33e98861a2400c4c42ed064cb82df097d41e5ff144dace786902e526fd2c67bb70ed91556d234d7d4902f13c936005d89d61086777546487b0f50cad1249e25ae7370ade106b52fa4f7eb3777fe841b9524bdafe9c39ce35e80ee39bdd9766b2cd5a7396d04a1d6e85ee034cb31a16e576a82515ad12eaa0a6a4b941da9ba3edfb8eb5fdc630ad87479fca12eafc14c6849e60001e2578ac6b1a0f8827eb9c0cdd15d6408c2778546cfebb66a3d86717c24448b9c28538ba063006b1801615f5a3;

endmodule

